module originalCU
(
	input CLOCK_50,
	input [9:0]SW, //SW[9] = sensor X
	input [1:0]KEY, //clock and clear
	output wire [9:0] LEDG, LEDR
);


parameter s0 = 3'b000, s1 = 3'b001, s2 = 3'b010, s3 = 3'b011, s4 = 3'b100;
parameter G = 2'b00, Y = 2'b01, R = 2'b10; 
reg [2:0]state, n_state;
reg [1:0]hwy, cntry;

assign LEDR [1:0] = hwy;
assign LEDG [1:0] = cntry;

assign LEDR [9:7] = state;

always@(negedge KEY[1], negedge KEY[0]) //clock and clear
	if(!KEY[0])
		state <= s0;
	else
		state <= n_state;
		

always@(state, SW[9])
begin
	case(state)
	s0: if(SW[9])
			n_state = s1;
		else
			n_state = s0;
	s1:	n_state = s2;
	s2: n_state = s3;
	s3: if(SW[9])
			n_state = s3;
		else
			n_state = s4;
	s4: n_state = s0;
	default: n_state = s0;
	endcase
end

always@(state)
begin
	case(state)
	s0: begin
		hwy = G;
		cntry = R;
		end
	s1: begin
		hwy = Y;
		cntry = R;
		end
	s2: begin
		hwy = R;
		cntry = R;
		end
	s3: begin
		hwy = R;
		cntry = G;
		end
	s4: begin
		hwy = R;
		cntry = Y;
		end
	endcase
end
endmodule

